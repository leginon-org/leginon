[x21] ; how many groups
; divides list into x21 evenly distributed groups
;  if x21=2 will divide into odd/even keys 
; retains only first register

FR
?IN.PARTICLE LIST TO DIVIDE (dir/doc)?<pcllist>
FR
?OUT.TEMPLATE FOR GROUP LISTS (dir/tmpl***)?<outtmpl>

; ~~~~~ start ~~~~~
UD N x22 ; number of particles
<pcllist>

VM
echo -n 'Dividing list of' {%F9.1%x22} 'particles into' {%F7.1%x21} 'groups..'

x30=x22 ; remaining particles
x40=0   ; particles processed
DO LB1 x11=1,x21  ; for each group

  x31=x30/(x21-x11+1) ;remaining particles / groups remaining
  x32=INT(x31) ;int(particles per group)
  x33=x31-x32  ;remainder

  IF(x33.gt.0)x32=x32+1 ;round up particles per group
  IF(x33.lt.0)THEN
    VM
    echo ERROR...negative remainder...END SCRIPT
    EN
  ENDIF

  SD IC NEW
  divpcllist_ic
  (1),x32 ;keys regs

  ;VM
  ;echo group {%F%x11} has {%F7.1%x32} particles
  DO LB2 x12=1,x32 ; for each particle in this group
    x34=x11+x21*(x12-1) ;key = group + interval * (round -1)

    UD IC x34,x35
    <pcllist>

    SD IC x12,x35
    divpcllist_ic

  LB2 ; next particle
  SD IC COPY
  divpcllist_ic
  <outtmpl>x11
  SD IC E
  divpcllist_ic

  x30=x30-x32 ; remaining particles

LB1
UD ICE
<pcllist>

VM
echo .done.

RE
